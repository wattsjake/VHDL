--standard library
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


entity full_adder is
  Port (X, Y, Cin: in std_logic;
		S, Co:     out std_logic);
end full_adder;

architecture Behavioral of full_adder is


begin



end Behavioral;
